module CoreTop(
    input clk
);












endmodule