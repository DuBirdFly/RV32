`include "defines.v"

module CoreTop(
    input clk
);












endmodule