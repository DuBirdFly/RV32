`include "defines.v"

module CoreTop(
    input                       clk,
    input                       rst
);

endmodule